module DrawEngine(input logic [31:0] AVL_READDATA,
	input logic [9:0] DrawY,
	output logic [9:0] AddrX, AddrY,
	output logic [15:0] ColorIdx,
	output logic [1:0] AVL_ADDR,			// Avalon-MM Address
	output logic [19:0] SRAM_ADDR,
	);
	

endmodule
